LavaStatus=0
   XM    �          j  e 
    j  e  T   
   ( �Gҡ��      o< 2       G         [ 2      ,2*   �   2         S h o o t e r . z i p m s e d g e . e x e h t t p s : / / d i g i l a b . d e i b . p o l i m i . i t / s / 8 c X a a 3 3 e k b s Q f p c / d o w n l o a d ? p a t h = % 2 F & f i l e s = S h o o t e r & d o w n l o a d S t a r t S e c r e t = 1 a 0 5 q g j g 8 s s (�R